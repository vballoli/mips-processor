module instruction_fetch()


endmodule